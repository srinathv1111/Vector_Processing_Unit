module Poly_Mul_Unit ();

endmodule